library verilog;
use verilog.vl_types.all;
entity sc_interrupt_vlg_vec_tst is
end sc_interrupt_vlg_vec_tst;
